package p1;
class c1;
int var1;
task t1(virtual mem_intf w1);
	var1=w1.rst;
endtask : t1
endclass
	
endpackage : p1